module sample_ploy_cbd;
endmodule