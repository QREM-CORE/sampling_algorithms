module sample_ntt;
endmodule