module tb_sample_poly_cbd;
endmodule