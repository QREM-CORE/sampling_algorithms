module tb_sample_ntt;
endmodule